typedef logic [31:0] word;
typedef logic [127:0] block;

